module Top_tb;

    Top dut();
    
    initial #800 $finish;
    

endmodule